* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_io__inv_1 A VGND VNB VPB VPWR Y
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1120000u l=150000u
.ends

.subckt sky130_fd_sc_io__nor2_1 A B VGND VNB VPB VPWR Y
X0 a_109_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1120000u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 Y B a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1120000u l=150000u
.ends

.subckt sky130_fd_sc_io__xor2_1 A B VGND VNB VPB VPWR X
X0 a_35_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND B a_35_297# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 X a_35_297# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_285_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1260000u l=150000u
X4 VPWR A a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1260000u l=150000u
X5 a_35_297# B a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1260000u l=150000u
X6 a_117_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1260000u l=150000u
X7 a_285_47# B X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_285_297# a_35_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1260000u l=150000u
X9 VGND A a_285_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends

.subckt sky130_fd_sc_io__nand2_1 A B VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1120000u l=150000u
X1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1120000u l=150000u
X2 VGND B a_113_47# VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
X3 a_113_47# A Y VNB sky130_fd_pr__nfet_01v8 w=740000u l=150000u
.ends

